module ScreenControl(wall_p1_xi, wall_p2_xi, LOC_p1_xi, LOC_p2_xi,wall_p1_yi, wall_p2_yi, LOC_p1_yi, LOC_p2_yi);
	parameter gridWidth = 8;
	parameter gridHeight = 8;
	input [gridWidth-1: 0] wall_p1_xi;
	input [gridWidth-1: 0] wall_p2_xi;
	input [gridWidth-1: 0] LOC_p1_xi;
	input [gridWidth-1: 0] LOC_p2_xi;
	input [gridHeight-1: 0] wall_p1_yi;
	input [gridHeight-1: 0] wall_p2_yi;
	input [gridHeight-1: 0] LOC_p1_yi;
	input [gridHeight-1: 0] LOC_p2_yi;
	
	

endmodule
