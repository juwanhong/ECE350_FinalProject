module Grid(enable1,enable2, clock, reset
,wall_p1_x, wall_p2_x, LOC_p1_x, LOC_p2_x,wall_p1_y, wall_p2_y, LOC_p1_y, LOC_p2_y
,wall_p1_xi, wall_p2_xi, LOC_p1_xi, LOC_p2_xi,wall_p1_yi, wall_p2_yi, LOC_p1_yi, LOC_p2_yi);
	parameter gridWidth = 32;
	parameter gridHeight = 32;
	input clock, enable1, enable2, reset;
	input [gridWidth-1: 0] wall_p1_xi;
	input [gridWidth-1: 0] wall_p2_xi;
	input [gridWidth-1: 0] LOC_p1_xi;
	input [gridWidth-1: 0] LOC_p2_xi;
	input [gridHeight-1: 0] wall_p1_yi;
	input [gridHeight-1: 0] wall_p2_yi;
	input [gridHeight-1: 0] LOC_p1_yi;
	input [gridHeight-1: 0] LOC_p2_yi;
	
	output [gridWidth-1: 0] wall_p1_x;
	output [gridWidth-1: 0] wall_p2_x;
	output [gridWidth-1: 0] LOC_p1_x;
	output [gridWidth-1: 0] LOC_p2_x;
	output [gridHeight-1: 0] wall_p1_y;
	output [gridHeight-1: 0] wall_p2_y;
	output [gridHeight-1: 0] LOC_p1_y;
	output [gridHeight-1: 0] LOC_p2_y;


genvar x,y;
generate
for (x = 0; x < gridWidth; x = x + 1)
begin: X
	DFFx df_x_p1_w(.d(wall_p1_xi[x]), .q(wall_p1_x[x]), .clk(clock), .en(enable1),.clrn(reset));
	DFFx df_x_p2_w(.d(wall_p2_xi[x]), .q(wall_p2_x[x]), .clk(clock), .en(enable2),.clrn(reset));
	DFFx df_x_p1_p(.d(LOC_p1_xi[x]), .q(LOC_p1_x[x]), .clk(clock), .en(enable1),.clrn(reset));
	DFFx df_x_p2_p(.d(LOC_p2_xi[x]), .q(LOC_p2_x[x]), .clk(clock), .en(enable2),.clrn(reset));

end
for (y = 0; y < gridHeight; y = y + 1)
begin: Y
	DFFx df_y_p1_w(.d(wall_p1_yi[y]), .q(wall_p1_y[y]), .clk(clock), .en(enable1),.clrn(reset));
	DFFx df_y_p2_w(.d(wall_p2_yi[y]), .q(wall_p2_y[y]), .clk(clock), .en(enable2),.clrn(reset));
	DFFx df_y_p1_p(.d(LOC_p1_yi[y]), .q(LOC_p1_y[y]), .clk(clock), .en(enable1),.clrn(reset));
	DFFx df_y_p2_p(.d(LOC_p2_yi[y]), .q(LOC_p2_y[y]), .clk(clock), .en(enable2),.clrn(reset));
end
endgenerate
endmodule

